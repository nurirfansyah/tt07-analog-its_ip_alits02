magic
tech sky130A
magscale 1 2
timestamp 1717269115
<< metal1 >>
rect 12080 12770 12440 12820
rect 12080 12540 12130 12770
rect 12390 12751 12440 12770
rect 12390 12609 18751 12751
rect 12390 12540 12440 12609
rect 12080 12490 12440 12540
rect 18613 12340 18747 12609
rect 18420 12280 18750 12340
rect 18050 12200 18750 12280
rect 18160 11940 19330 12040
rect 19232 11620 19328 11940
rect 19140 11580 19400 11620
rect 19140 11400 19180 11580
rect 19360 11400 19400 11580
rect 19140 11370 19400 11400
rect 17880 9126 18100 9140
rect 14664 8926 14670 9126
rect 14870 8926 15310 9126
rect 17880 8926 17892 9126
rect 18092 8926 18100 9126
rect 17880 8910 18100 8926
rect 16110 6610 16420 7910
rect 17000 7300 17280 7900
rect 17000 7240 17360 7300
rect 17000 7010 17060 7240
rect 17300 7010 17360 7240
rect 17000 6970 17360 7010
rect 16110 6390 16160 6610
rect 16370 6390 16420 6610
rect 16110 6350 16420 6390
rect 14664 5510 14670 5710
rect 14870 5510 14876 5710
rect 20354 5510 20360 5710
rect 20560 5510 20566 5710
rect 14670 1560 14870 5510
rect 20360 2250 20560 5510
rect 21830 5100 23190 5130
rect 28100 5110 29480 5190
rect 21830 4990 21880 5100
rect 23140 5080 23190 5100
rect 23140 5000 28310 5080
rect 23140 4990 23190 5000
rect 21830 4960 23190 4990
rect 28780 4840 28930 4860
rect 28600 4740 28800 4840
rect 28900 4740 28930 4840
rect 28780 4710 28930 4740
rect 29310 4600 29480 5110
rect 25130 4490 25340 4520
rect 25130 4400 25150 4490
rect 25310 4480 25340 4490
rect 25310 4400 25900 4480
rect 29310 4460 29330 4600
rect 29460 4460 29480 4600
rect 29310 4440 29480 4460
rect 25130 4380 25340 4400
rect 20360 2044 20560 2050
rect 14670 1360 27840 1560
rect 27640 1090 27840 1360
rect 27550 1030 27930 1090
rect 27550 760 27610 1030
rect 27870 760 27930 1030
rect 27550 710 27930 760
<< via1 >>
rect 12130 12540 12390 12770
rect 19180 11400 19360 11580
rect 14670 8926 14870 9126
rect 17892 8926 18092 9126
rect 17060 7010 17300 7240
rect 16160 6390 16370 6610
rect 14670 5510 14870 5710
rect 20360 5510 20560 5710
rect 21880 4990 23140 5100
rect 28800 4740 28900 4840
rect 25150 4400 25310 4490
rect 29330 4460 29460 4600
rect 20360 2050 20560 2250
rect 27610 760 27870 1030
<< metal2 >>
rect 50 12770 12440 12820
rect 50 12760 12130 12770
rect 50 12540 140 12760
rect 550 12540 12130 12760
rect 12390 12540 12440 12770
rect 50 12490 12440 12540
rect 19140 11580 19400 11620
rect 19140 11400 19180 11580
rect 19360 11400 19400 11580
rect 19140 11370 19400 11400
rect 14670 9126 14870 9132
rect 14670 5710 14870 8926
rect 17880 9126 18100 9140
rect 17880 8926 17892 9126
rect 18092 8926 20560 9126
rect 17880 8910 18100 8926
rect 17000 7240 17360 7300
rect 17000 7010 17060 7240
rect 17300 7010 17360 7240
rect 17000 6970 17360 7010
rect 16110 6610 16420 6670
rect 16110 6390 16160 6610
rect 16370 6390 16420 6610
rect 16110 6350 16420 6390
rect 14670 5504 14870 5510
rect 20360 5710 20560 8926
rect 20360 5504 20560 5510
rect 140 5150 23230 5190
rect 140 4820 170 5150
rect 500 5100 23230 5150
rect 500 4990 21880 5100
rect 23140 4990 23230 5100
rect 500 4820 23230 4990
rect 140 4790 23230 4820
rect 28780 4850 31490 4870
rect 28780 4840 31280 4850
rect 28780 4740 28800 4840
rect 28900 4740 31280 4840
rect 28780 4730 31280 4740
rect 31440 4730 31490 4850
rect 28780 4710 31490 4730
rect 29290 4600 29500 4620
rect 25130 4490 25340 4520
rect 25130 4400 25150 4490
rect 25310 4400 25340 4490
rect 29290 4460 29330 4600
rect 29460 4460 29500 4600
rect 29290 4440 29500 4460
rect 25130 4380 25340 4400
rect 9710 3720 28630 3770
rect 9710 3250 9760 3720
rect 10140 3250 28630 3720
rect 9710 3190 28630 3250
rect 20354 2050 20360 2250
rect 20560 2050 20566 2250
rect 20360 1010 20560 2050
rect 22410 1030 25330 1050
rect 27550 1030 27930 1090
rect 22410 1010 22460 1030
rect 20360 850 22460 1010
rect 22640 850 25160 1030
rect 25290 850 25330 1030
rect 20360 830 25330 850
rect 26790 1010 27610 1030
rect 26790 840 26860 1010
rect 27040 840 27610 1010
rect 20360 810 22990 830
rect 26790 820 27610 840
rect 27550 760 27610 820
rect 27870 1010 29550 1030
rect 27870 840 29320 1010
rect 29500 840 29550 1010
rect 27870 820 29550 840
rect 27870 760 27930 820
rect 27550 710 27930 760
<< via2 >>
rect 140 12540 550 12760
rect 19180 11400 19360 11580
rect 17060 7010 17300 7240
rect 16160 6390 16370 6610
rect 170 4820 500 5150
rect 31280 4730 31440 4850
rect 25150 4400 25310 4490
rect 29330 4460 29460 4600
rect 9760 3250 10140 3720
rect 22460 850 22640 1030
rect 25160 850 25290 1030
rect 26860 840 27040 1010
rect 29320 840 29500 1010
<< metal3 >>
rect 80 12760 610 12820
rect 80 12540 140 12760
rect 550 12540 610 12760
rect 80 12490 610 12540
rect 19095 11580 19425 11665
rect 19095 11400 19180 11580
rect 19360 11400 19425 11580
rect 17000 7240 17360 7300
rect 17000 7010 17060 7240
rect 17300 7010 17360 7240
rect 17000 6970 17360 7010
rect 17930 6975 18340 7020
rect 19095 6975 19425 11400
rect 16110 6610 16420 6670
rect 16110 6390 16160 6610
rect 16370 6390 16420 6610
rect 16110 6350 16420 6390
rect 17930 6645 19425 6975
rect 140 5150 540 5190
rect 140 4820 170 5150
rect 500 4820 540 5150
rect 140 4790 540 4820
rect 9710 3720 10200 3770
rect 9710 3250 9760 3720
rect 10140 3250 10200 3720
rect 9710 3190 10200 3250
rect 17930 2870 18260 6645
rect 31260 4850 31460 4890
rect 31260 4730 31280 4850
rect 31440 4730 31460 4850
rect 29310 4600 29480 4620
rect 25140 4520 25310 4560
rect 25130 4490 25340 4520
rect 25130 4400 25150 4490
rect 25310 4400 25340 4490
rect 25130 4380 25340 4400
rect 29310 4460 29330 4600
rect 29460 4460 29480 4600
rect 17930 2300 18020 2870
rect 18190 2300 18260 2870
rect 17930 2280 18260 2300
rect 22440 1030 22660 1100
rect 22440 850 22460 1030
rect 22640 850 22660 1030
rect 22440 470 22660 850
rect 25140 1030 25310 4380
rect 25140 850 25160 1030
rect 25290 850 25310 1030
rect 25140 830 25310 850
rect 26840 1010 27060 1060
rect 29310 1030 29480 4460
rect 26840 840 26860 1010
rect 27040 840 27060 1010
rect 22420 450 22670 470
rect 22420 310 22440 450
rect 22650 310 22670 450
rect 22420 290 22670 310
rect 26840 440 27060 840
rect 29300 1010 29520 1030
rect 29300 840 29320 1010
rect 29500 840 29520 1010
rect 29300 820 29520 840
rect 31260 440 31460 4730
rect 26840 420 27080 440
rect 26840 310 26860 420
rect 27050 310 27080 420
rect 26840 290 27080 310
rect 31260 310 31280 440
rect 31440 310 31460 440
rect 31260 290 31460 310
<< via3 >>
rect 140 12540 550 12760
rect 17060 7010 17300 7240
rect 16160 6390 16370 6610
rect 170 4820 500 5150
rect 9760 3250 10140 3720
rect 18020 2300 18190 2870
rect 22440 310 22650 450
rect 26860 310 27050 420
rect 31280 310 31440 440
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 760 44820 11948 44952
rect 200 12820 500 44152
rect 80 12760 610 12820
rect 80 12540 140 12760
rect 550 12540 610 12760
rect 80 12490 610 12540
rect 200 5190 500 12490
rect 9800 10800 10100 44820
rect 9800 10510 16480 10800
rect 140 5150 540 5190
rect 140 4820 170 5150
rect 500 4820 540 5150
rect 140 4790 540 4820
rect 200 1000 500 4790
rect 9800 3770 10100 10510
rect 17000 7240 17360 7300
rect 17000 7010 17060 7240
rect 17300 7010 17360 7240
rect 17000 6970 17360 7010
rect 16110 6610 16420 6670
rect 16110 6390 16160 6610
rect 16370 6390 16420 6610
rect 16110 6350 16420 6390
rect 16205 4225 16415 6350
rect 12415 4015 16415 4225
rect 9710 3720 10200 3770
rect 9710 3250 9760 3720
rect 10140 3250 10200 3720
rect 9710 3190 10200 3250
rect 9800 1000 10100 3190
rect 12415 410 12625 4015
rect 13595 2704 13805 2705
rect 17044 2704 17254 6970
rect 13595 2497 17254 2704
rect 13595 410 13805 2497
rect 17044 2495 17254 2497
rect 18001 2870 18209 2894
rect 18001 2300 18020 2870
rect 18190 2300 18209 2870
rect 18001 410 18209 2300
rect 22420 450 22670 470
rect 9150 200 12635 410
rect 13580 200 13840 410
rect 18000 200 18260 410
rect 22420 310 22440 450
rect 22650 310 22670 450
rect 31260 440 31490 460
rect 22420 290 22670 310
rect 26840 420 27070 440
rect 26840 310 26860 420
rect 27050 310 27070 420
rect 26840 290 27070 310
rect 31260 310 31280 440
rect 31440 310 31490 440
rect 31260 290 31490 310
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 290
rect 26866 0 27046 290
rect 31282 0 31462 290
use pll  pll_0 ~/design/irfan/tt07-analog-its_ip_alits02/mag/dsrt_pll
timestamp 1717268110
transform 1 0 14390 0 1 9446
box -230 -1596 4416 5184
use vco  vco_0 ~/design/irfan/tt07-analog-its_ip_alits02/mag/dsrt_vco
timestamp 1717263762
transform 1 0 25450 0 1 3880
box -600 -1710 3900 3550
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
