magic
tech sky130A
timestamp 1717262129
<< metal1 >>
rect 14655 2595 14735 2615
rect 10915 2550 11595 2565
rect 14050 2555 14665 2595
rect 10915 2495 10940 2550
rect 11570 2540 11595 2550
rect 14655 2545 14665 2555
rect 14725 2545 14735 2595
rect 11570 2500 14155 2540
rect 14655 2535 14735 2545
rect 11570 2495 11595 2500
rect 10915 2480 11595 2495
rect 14390 2420 14465 2430
rect 14300 2370 14400 2420
rect 14450 2370 14465 2420
rect 14390 2355 14465 2370
rect 12565 2245 12670 2260
rect 12565 2200 12575 2245
rect 12655 2240 12670 2245
rect 12655 2200 12950 2240
rect 12565 2190 12670 2200
<< via1 >>
rect 10940 2495 11570 2550
rect 14665 2545 14725 2595
rect 14400 2370 14450 2420
rect 12575 2200 12655 2245
<< metal2 >>
rect 14655 2595 14735 2615
rect 70 2575 11615 2595
rect 70 2410 85 2575
rect 250 2550 11615 2575
rect 250 2495 10940 2550
rect 11570 2495 11615 2550
rect 14655 2535 14665 2595
rect 14725 2535 14735 2595
rect 14655 2525 14735 2535
rect 250 2410 11615 2495
rect 70 2395 11615 2410
rect 14390 2425 15745 2435
rect 14390 2420 15640 2425
rect 14390 2370 14400 2420
rect 14450 2370 15640 2420
rect 14390 2365 15640 2370
rect 15720 2365 15745 2425
rect 14390 2355 15745 2365
rect 12565 2245 12670 2260
rect 12565 2200 12575 2245
rect 12655 2200 12670 2245
rect 12565 2190 12670 2200
rect 4855 1860 14315 1885
rect 4855 1625 4880 1860
rect 5070 1625 14315 1860
rect 4855 1595 14315 1625
rect 11205 515 12665 525
rect 11205 425 11230 515
rect 11320 425 12580 515
rect 12645 425 12665 515
rect 11205 415 12665 425
rect 13395 505 14775 515
rect 13395 420 13430 505
rect 13520 420 14660 505
rect 14750 420 14775 505
rect 13395 410 14775 420
<< via2 >>
rect 85 2410 250 2575
rect 14665 2545 14725 2585
rect 14665 2535 14725 2545
rect 15640 2365 15720 2425
rect 12575 2200 12655 2245
rect 4880 1625 5070 1860
rect 11230 425 11320 515
rect 12580 425 12645 515
rect 13430 420 13520 505
rect 14660 420 14750 505
<< metal3 >>
rect 70 2575 270 2595
rect 70 2410 85 2575
rect 250 2410 270 2575
rect 70 2395 270 2410
rect 14655 2585 14740 2595
rect 14655 2535 14665 2585
rect 14725 2535 14740 2585
rect 12570 2260 12655 2280
rect 12565 2245 12670 2260
rect 12565 2200 12575 2245
rect 12655 2200 12670 2245
rect 12565 2190 12670 2200
rect 4855 1860 5100 1885
rect 4855 1625 4880 1860
rect 5070 1625 5100 1860
rect 4855 1595 5100 1625
rect 11220 515 11330 550
rect 11220 425 11230 515
rect 11320 425 11330 515
rect 11220 235 11330 425
rect 12570 515 12655 2190
rect 12570 425 12580 515
rect 12645 425 12655 515
rect 12570 415 12655 425
rect 13420 505 13530 530
rect 14655 515 14740 2535
rect 15630 2425 15730 2445
rect 15630 2365 15640 2425
rect 15720 2365 15730 2425
rect 13420 420 13430 505
rect 13520 420 13530 505
rect 11210 225 11335 235
rect 11210 155 11220 225
rect 11325 155 11335 225
rect 11210 145 11335 155
rect 13420 220 13530 420
rect 14650 505 14760 515
rect 14650 420 14660 505
rect 14750 420 14760 505
rect 14650 410 14760 420
rect 15630 220 15730 2365
rect 13420 210 13540 220
rect 13420 155 13430 210
rect 13525 155 13540 210
rect 13420 145 13540 155
rect 15630 155 15640 220
rect 15720 155 15730 220
rect 15630 145 15730 155
<< via3 >>
rect 85 2410 250 2575
rect 4880 1625 5070 1860
rect 11220 155 11325 225
rect 13430 155 13525 210
rect 15640 155 15720 220
<< metal4 >>
rect 399 22476 429 22576
rect 767 22476 797 22576
rect 1135 22476 1165 22576
rect 1503 22476 1533 22576
rect 1871 22476 1901 22576
rect 2239 22476 2269 22576
rect 2607 22476 2637 22576
rect 2975 22476 3005 22576
rect 3343 22476 3373 22576
rect 3711 22476 3741 22576
rect 4079 22476 4109 22576
rect 4447 22476 4477 22576
rect 4815 22476 4845 22576
rect 5183 22476 5213 22576
rect 5551 22476 5581 22576
rect 5919 22476 5949 22576
rect 6287 22476 6317 22576
rect 6655 22476 6685 22576
rect 7023 22476 7053 22576
rect 7391 22476 7421 22576
rect 7759 22476 7789 22576
rect 8127 22476 8157 22576
rect 8495 22476 8525 22576
rect 8863 22476 8893 22576
rect 9231 22476 9261 22576
rect 9599 22476 9629 22576
rect 9967 22476 9997 22576
rect 10335 22476 10365 22576
rect 10703 22476 10733 22576
rect 11071 22476 11101 22576
rect 11439 22476 11469 22576
rect 11807 22476 11837 22576
rect 12175 22476 12205 22576
rect 12543 22476 12573 22576
rect 12911 22476 12941 22576
rect 13279 22476 13309 22576
rect 13647 22476 13677 22576
rect 14015 22476 14045 22576
rect 14383 22476 14413 22576
rect 14751 22476 14781 22576
rect 15119 22476 15149 22576
rect 15487 22476 15517 22576
rect 15855 22476 15885 22576
rect 100 2595 250 22076
rect 70 2575 270 2595
rect 70 2410 85 2575
rect 250 2410 270 2575
rect 70 2395 270 2410
rect 100 500 250 2395
rect 4900 1885 5050 22076
rect 4855 1860 5100 1885
rect 4855 1625 4880 1860
rect 5070 1625 5100 1860
rect 4855 1595 5100 1625
rect 4900 500 5050 1595
rect 11210 225 11335 235
rect 11210 155 11220 225
rect 11325 155 11335 225
rect 15630 220 15745 230
rect 11210 145 11335 155
rect 13420 210 13535 220
rect 13420 155 13430 210
rect 13525 155 13535 210
rect 13420 145 13535 155
rect 15630 155 15640 220
rect 15720 155 15745 220
rect 15630 145 15745 155
rect 185 0 275 100
rect 2393 0 2483 100
rect 4601 0 4691 100
rect 6809 0 6899 100
rect 9017 0 9107 100
rect 11225 0 11315 145
rect 13433 0 13523 145
rect 15641 0 15731 145
use vco  vco_0 ~/design/irfan/tt07-analog-its_ip_alits02/mag/dsrt_vco
timestamp 1717229036
transform 1 0 12725 0 1 1940
box -300 -855 1950 1775
<< labels >>
flabel metal4 s 15487 22476 15517 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 15855 22476 15885 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 15119 22476 15149 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15641 0 15731 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13433 0 13523 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11225 0 11315 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9017 0 9107 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 6809 0 6899 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 4601 0 4691 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 2393 0 2483 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 185 0 275 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 14751 22476 14781 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 14015 22476 14045 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13647 22476 13677 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12911 22476 12941 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12543 22476 12573 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11807 22476 11837 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11439 22476 11469 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10703 22476 10733 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10335 22476 10365 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9599 22476 9629 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9231 22476 9261 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 2975 22476 3005 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 2607 22476 2637 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 2239 22476 2269 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 1871 22476 1901 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 1503 22476 1533 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 1135 22476 1165 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 767 22476 797 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 399 22476 429 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 5919 22476 5949 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 5183 22476 5213 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 4815 22476 4845 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 4079 22476 4109 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 3711 22476 3741 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 8495 22476 8525 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8127 22476 8157 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 7391 22476 7421 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 7023 22476 7053 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 6287 22476 6317 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 250 22076 1 FreeSans 1 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 4900 500 5050 22076 1 FreeSans 1 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
