VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_nurirfansyah_alits02
  CLASS BLOCK ;
  FOREIGN tt_um_nurirfansyah_alits02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.810000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 127.850 24.000 129.350 25.650 ;
        RECT 130.650 24.000 132.150 25.650 ;
        RECT 133.450 24.000 134.950 25.650 ;
        RECT 136.250 24.000 137.750 25.650 ;
        RECT 139.050 24.000 140.550 25.650 ;
        RECT 141.850 24.000 143.350 25.650 ;
      LAYER li1 ;
        RECT 128.050 25.100 128.600 25.400 ;
        RECT 128.800 25.000 129.350 25.950 ;
        RECT 130.850 25.100 131.950 25.400 ;
        RECT 133.650 25.100 134.200 25.400 ;
        RECT 128.050 23.200 128.450 24.850 ;
        RECT 128.750 24.150 129.150 24.750 ;
        RECT 130.850 24.300 131.250 25.100 ;
        RECT 133.650 25.000 134.050 25.100 ;
        RECT 134.400 25.000 134.950 25.950 ;
        RECT 136.450 25.100 137.550 25.400 ;
        RECT 139.250 25.100 139.800 25.400 ;
        RECT 128.750 23.750 129.350 24.150 ;
        RECT 130.650 23.850 131.300 24.100 ;
        RECT 128.750 23.200 129.150 23.750 ;
        RECT 128.050 22.550 128.600 22.850 ;
        RECT 128.800 22.000 129.350 22.950 ;
        RECT 130.850 22.850 131.250 23.650 ;
        RECT 131.550 23.200 131.950 24.750 ;
        RECT 133.650 23.200 134.050 24.750 ;
        RECT 134.350 24.150 134.750 24.750 ;
        RECT 136.450 24.300 136.850 25.100 ;
        RECT 139.250 25.000 139.650 25.100 ;
        RECT 140.000 25.000 140.550 25.950 ;
        RECT 142.050 25.100 143.150 25.400 ;
        RECT 134.350 23.750 134.950 24.150 ;
        RECT 136.250 23.850 136.900 24.100 ;
        RECT 134.350 23.200 134.750 23.750 ;
        RECT 130.850 22.550 131.950 22.850 ;
        RECT 133.650 22.550 134.200 22.850 ;
        RECT 134.400 22.000 134.950 22.950 ;
        RECT 136.450 22.850 136.850 23.650 ;
        RECT 137.150 23.200 137.550 24.750 ;
        RECT 139.250 23.200 139.650 24.750 ;
        RECT 139.950 24.150 140.350 24.750 ;
        RECT 142.050 24.300 142.450 25.100 ;
        RECT 139.950 23.750 140.550 24.150 ;
        RECT 141.850 23.850 142.500 24.100 ;
        RECT 139.950 23.200 140.350 23.750 ;
        RECT 136.450 22.550 137.550 22.850 ;
        RECT 139.250 22.550 139.800 22.850 ;
        RECT 140.000 22.000 140.550 22.950 ;
        RECT 142.050 22.850 142.450 23.650 ;
        RECT 142.750 23.200 143.150 24.750 ;
        RECT 142.050 22.550 143.150 22.850 ;
      LAYER met1 ;
        RECT 146.550 25.950 147.350 26.150 ;
        RECT 109.150 25.400 115.950 25.650 ;
        RECT 128.050 25.550 147.350 25.950 ;
        RECT 109.150 25.000 143.150 25.400 ;
        RECT 146.550 25.350 147.350 25.550 ;
        RECT 109.150 24.800 115.950 25.000 ;
        RECT 128.050 24.350 143.150 24.750 ;
        RECT 128.050 23.600 128.450 24.350 ;
        RECT 142.750 24.200 143.150 24.350 ;
        RECT 143.900 24.200 144.650 24.300 ;
        RECT 128.750 23.750 131.300 24.200 ;
        RECT 131.550 23.750 134.050 24.200 ;
        RECT 134.350 23.750 136.900 24.200 ;
        RECT 137.150 23.750 139.650 24.200 ;
        RECT 139.950 23.750 142.500 24.200 ;
        RECT 142.750 23.700 144.650 24.200 ;
        RECT 142.750 23.600 143.150 23.700 ;
        RECT 128.050 23.200 143.150 23.600 ;
        RECT 143.900 23.550 144.650 23.700 ;
        RECT 125.650 22.400 126.700 22.600 ;
        RECT 128.050 22.550 143.150 22.950 ;
        RECT 125.650 22.000 140.550 22.400 ;
        RECT 125.650 21.900 126.700 22.000 ;
        RECT 140.750 15.950 143.150 22.550 ;
      LAYER met2 ;
        RECT 0.700 23.950 116.150 25.950 ;
        RECT 146.550 25.250 147.350 26.150 ;
        RECT 129.250 23.750 130.750 24.200 ;
        RECT 134.850 23.750 136.350 24.200 ;
        RECT 140.450 23.750 141.950 24.200 ;
        RECT 143.900 23.550 157.450 24.350 ;
        RECT 125.650 21.900 126.700 22.600 ;
        RECT 140.750 18.850 143.150 21.050 ;
        RECT 48.550 15.950 143.150 18.850 ;
        RECT 112.050 4.150 126.650 5.250 ;
        RECT 133.950 4.100 147.750 5.150 ;
      LAYER met3 ;
        RECT 124.250 26.650 134.700 37.100 ;
        RECT 136.300 26.700 146.750 37.150 ;
        RECT 0.700 23.950 2.700 25.950 ;
        RECT 129.250 23.750 130.750 26.650 ;
        RECT 125.700 22.600 126.550 22.800 ;
        RECT 125.650 21.900 126.700 22.600 ;
        RECT 48.550 15.950 51.000 18.850 ;
        RECT 112.200 2.350 113.300 5.500 ;
        RECT 125.700 4.150 126.550 21.900 ;
        RECT 134.850 21.250 136.350 24.200 ;
        RECT 140.450 23.750 141.950 26.700 ;
        RECT 129.650 10.850 140.050 21.250 ;
        RECT 140.750 15.950 143.150 21.050 ;
        RECT 112.100 1.450 113.350 2.350 ;
        RECT 134.200 2.200 135.300 5.300 ;
        RECT 146.550 5.150 147.400 25.950 ;
        RECT 146.500 4.100 147.600 5.150 ;
        RECT 134.200 1.450 135.400 2.200 ;
        RECT 156.300 1.450 157.300 24.450 ;
      LAYER met4 ;
        RECT 124.600 31.500 129.350 31.550 ;
        RECT 124.600 27.000 146.500 31.500 ;
        RECT 124.600 26.950 129.350 27.000 ;
        RECT 0.700 23.950 1.000 25.950 ;
        RECT 2.500 23.950 2.700 25.950 ;
        RECT 134.700 21.050 139.700 27.000 ;
        RECT 48.550 15.950 49.000 18.850 ;
        RECT 50.500 15.950 51.000 18.850 ;
        RECT 134.650 15.950 143.150 21.050 ;
        RECT 134.650 15.900 139.850 15.950 ;
        RECT 112.100 1.450 113.350 2.350 ;
        RECT 134.200 1.450 135.350 2.200 ;
        RECT 156.300 1.450 157.450 2.300 ;
        RECT 112.250 1.000 113.150 1.450 ;
        RECT 134.330 1.000 135.230 1.450 ;
        RECT 156.410 1.000 157.310 1.450 ;
  END
END tt_um_nurirfansyah_alits02
END LIBRARY

